�PNG

   IHDR           szz�  �IDATx�c|d	��b�<۶m۶m�6µm{c۶���훳��Pɠ����ɿU�8�	�p8� N�O�-?�I�X^L�Z'�[,S,���hH�X��c��{�s��$`�? N�XnV�©aam��7Xr��*6�r[-w��:�/9�,�y$���Д���dèS�)@���4��||�3�>��I�:�}��j�t�l<�D6}4�=�5����ߟU�ʃf�i��䨣�r�m�yx�hK�4��/��J5���������l��֌�bV�/kԠt�=����\ٿ(,�w}B���d��X��,eAL�Wv�q\���I@�'�v?	�9�y��֘w�)���Β�b~~,V�=�����^m�]U��F�-]��'鳢$����ՙ���pntqa�������F�nS�?
�
��8����s�aN@ 3�ܘ��m�a��֞��>��c�|�'w	�mMX���r���,//��+7�;U#�D�0�ǧ���ؤ����yZcFT�zzv}�¿��jr��������v�el��"��Kd�����G} x����G:����g�G�P7��
&�I��sR�����7ʌ�'�̆c�e�>�0O'��e
p�� tө�"�i��W���,ww�uu���H%a����7���7?Wl���h��ƲB^(��4D�Κ�At?XH�T��\++��d.Q�t�LW��r�6x>�K�6��M��y}t���f)wFD�	`�|�N�h�c�! V���*ꖅ2�̭��\%��������[�� 0�x: ~@^�^�UN���7�ͭ{��;:L|<�)0�� �7��R=<zS�V5D�{��G�'��+�� .�\D.f\�I���q�;��π�d��g��W��Z�Oru X$�G�������0F��¥@s:�/������0)J��8\�?)q�)=$�%[�6ǝ$�7=��C��Q�c'��%��/*	    IEND�B`�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           <svg xmlns="http://www.w3.org/2000/svg" width="22" height="22" version="1">
 <path style="opacity:0.05" d="m 2,1.5 c -0.554,0 -1,0.446 -1,1 V 11 H 21 V 2.5 c 0,-0.554 -0.446,-1 -1,-1 z"/>
 <rect style="fill:#687df9" width="20" height="20" x="1" y="1" rx="1" ry="1"/>
 <path style="opacity:0.2" d="M 9.8571,18.5 C 9.5406,18.5 8.9899,18.2597 9,17.9615 V 9.5 H 7 l 4,-5 4,5 h -2 v 8.4615 C 13,18.2598 12.459,18.5 12.143,18.5 Z"/>
 <path style="fill:#ffffff" d="M 9.8571,18 C 9.5406,18 8.9899,17.7597 9,17.4615 V 9 H 7 l 4,-5 4,5 h -2 v 8.4615 C 13,17.7598 12.459,18 12.143,18 Z"/>
 <path style="opacity:0.2;fill:#ffffff" d="M 1,2.5 V 2 C 1,1.446 1.446,1 2,1 h 18 c 0.554,0 1,0.446 1,1 v 0.5 c 0,-0.554 -0.446,-1 -1,-1 H 2 c -0.554,0 -1,0.446 -1,1 z"/>
 <path style="opacity:0.2" d="m 1,20 v 0.5 c 0,0.554 0.446,1 1,1 h 18 c 0.554,0 1,-0.446 1,-1 V 20 c 0,0.554 -0.446,1 -1,1 H 2 C 1.446,21 1,20.554 1,20 Z"/>
</svg>
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               <svg xmlns="http://www.w3.org/2000/svg" width="24" height="24" version="1.1">
 <defs>
  <style id="current-color-scheme" type="text/css">
   .ColorScheme-Text { color:#ffffff; } .ColorScheme-Highlight { color:#4285f4; } .ColorScheme-NeutralText { color:#ff9800; } .ColorScheme-PositiveText { color:#4caf50; } .ColorScheme-NegativeText { color:#f44336; }
  </style>
 </defs>
 <g style="fill:currentColor" class="ColorScheme-Text" transform="translate(3,-1029.4)">
  <rect width="8" height="15" x="5" y="1034.4" rx="1" ry="1"/>
  <path d="m2.25 1035.4c-0.1385 0-0.25 0.1115-0.25 0.25v0.5c0 0.1385 0.1115 0.25 0.25 0.25h1.75v-1h-1.75zm0 2c-0.1385 0-0.25 0.1115-0.25 0.25v0.5c0 0.1385 0.1115 0.25 0.25 0.25h1.75v-1h-1.75zm0 2c-0.1385 0-0.25 0.1115-0.25 0.25v0.5c0 0.1385 0.1115 0.25 0.25 0.25h1.75v-1h-1.7