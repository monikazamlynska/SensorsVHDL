A��!Y����u��Y�(c���r������*�y+)��b�S��O�}2�q@a�H'��&��q�˛���"����N��!g�B�(z$���J�	���u}�!˿>��!��0�������s !)�����'Յa�ro���>Qݬ��q��k�]��E�}�V��#[2�^�/�+��?J�-)�LU1�da��E¦�4���5s����U���E����E�����[�jt,���XܭvKM �� �3T�.�>/}?X��rdpf����cc�Sq[k�PL�m7=������>�vmF|�]����6��z(�����ae1�O�W�M<C6�ꄚZ
)�
��+�?�c-Y��ͷ��f���+h�P�ɽ���҅�b���5Y*��Fr�U��� io��`��oA���b�F���m�J�hz��҅���_��bs)ܻ¥jb�-��-p#c��{�pʒ�eU��Z���Q����
�d� ��#�q�[r�[��P��n�`?����~~��T��l��U���9a�Li�i�"�s-��>�A� ޤ
%�b�%d�$�	ҐV8�ĉ"
�y��T���e��y���0���A<ۧwm�l��_H��ۧ�.�?���R`1xX��1�o
ʎ���ە(]M�V�l���M�]!�[�#��z��g���V��ۉ�m�f�*��N�̅[8��M�d)m�d�%.���669�ff�M3;���.�{_Z�iQxvrh׾��z nW/��:�L�M'�6�ehZ�'�id���B�����rS��&;��`�<���	�;(��UN,8m��T�3�������G�m�}�-lu�ʠ|�J^WXn��AV�דWE���'7Ӑ[����4�k/t�J��#�M��9�Mv,kF�eE����ڂ�ŝRBY]2JY��`_+( ���WQxN��ɢ�C�kQ��R�Q��II�e���q>*����+b�-��v���U
!��������l[�ƙ匂$�b�j1��&�u���ʽ*�.c����7b��Gf��]�7tۥ���l�Ѧ���� 10��W�|�JZҦ�J���!ټn�ְ�h�� Nq����V��z�0u;1ZZ"@�Y�w�5���5�{Y��yU���>�{�h�,���Z[��m�3o��V)Z�>��ZtmZ�vtD��o�#`�� pIj�*䗄�<-U����92v[|.*� ��[@8+E~�fM��hF;K��9��ط���� @�q����b�YO�R$��s.���3&��v�v�������
6�S݌��).ⶋu/Ҭ=c�دMcL�J9��M.3�|3��!�q>w!���v�/��__��_-3!٫M�Y(�4!��U��#a����!��<TU\�t4��cD���q���2o��\���@8�w�aqg��R��,��gl�q�M��Zg�^r�5�͘hY%�%[�&��fSI��Ք�Ub���Hz�lI���i�k�Y_����yOH]�)�=s���6k�6�B]'q|n��i�X>hj�?�m�����/c��t:��?�r=|�ů�6 $�7�?(�/	�!�������ב���n���^��ns|ye[E�������w X�K��rx��U�5�.vTP,��)K����e�^|�F	.�=�t��zf����ړ��5z����L��cA�ƶh�[U`SK�]%�w�%�}<H� �g�;�mps��K��9�!��
L��j�Kğ}��v��H��M ��j�y��"�2�1��cw�G�d�)x�?�6�����!���QWK�Tß��+tu�#okf���"���3}�٘f��� ���Ow	��$�HK�m�}a�ش�r꺚�;���en4Ń�;�滍G1��5�|���Newm&�x�i�,��h\�����t�WW �0��\.�W�;�XE��>�~Ba3��1�7����B|߇p8p�q<��Jp0�@�L+8�#�
0�`!0f �b���P���4���<�����>�:R:�p����V�trA��<Y{�S�>�a�� ���� ���ڈ7�ߣdl��,1nU}�2P��X"�X��Ui�=� wg�y�b	�~	��	�r�[V�s�C���Ʌ�V���F����M�9Dv��ş����?�L��J��w�aAշ�
�`B��X�7�O�&>s�0uz=�u.}y���}m`Ң*%.׬��|�%2��F���e�1o,��	���a�+`A�/�1���^�@�L�<C�ż�5ʻ�d��H�f�
�z��o�B�rm4Vmj�(�j,uG�/m�Y�q��DB?Y�����QӃZ{ȃ�	Ё�!鼨*���G��&K6�ڛ~4�����C��h�G�1W=
m���[������n��'�I����gd�dȓ�1�s����{~�m~~ J�;���)�6���z�_%U��=�뻥� ��лi��%A�]��������U^�Nd�~��A]z��n�����ڀg��H����i.c���_�ձ.�+]W�U,ǝA���{����|�1ƿ �ۂH?=S��@e'��I>&L����>�c�(:=<��|š�DZB�c'vAߨ��W(�w�k �g�ܮ��ΫՅ~Wx���VO�|��j��۳�k���e�沛��db?�������e�	�r��j$���t�\�FtJ�Z�����?r9���6�����2D�,�eK+GS�Ԏ��/���g�{�!�rp� r��b��y���_��������vpဃ�r�.-Z�-������X����D�{�bw��b� �2-�6��ph۠�i�I�����5Bl�H���&�B �����<���=X�t�[z�t��󽌉�HC.��υ�~�ه�>o��>��}<��g� /��+�#_W	���q���޾N�Dz�I�衜>���up쟼�ט���e6�z��+Γ���	��$�����{�5���jq͓���\��h�z��ˇsr.�����ݤ���Y3��pC3��S{t�C��v���qp�~�N�����|-p�=����(gqd��~vrL � �g��E`�Y�1,�0�VHۈ�O��D���=�2�v�i��42[���M!/�w�5��7�
@�MDmM^���՛e��o�	���O��%)>��}DQ�	ٞ
�;Vu@�>,|nځk~��՝1GP(F��I�W�f���������Xu���i�&���A[�������ęI�����}0��%��5Cf&��̙\$_u9H�5��5�[�9v$��#�����$]�����p<^�肸�{�8��2����}yG�~n������KȺS	��o�ChvyV� ̠�.��JA���1���e���ʊ��x��� �p�B�İ$�a�0�a {#�&���N�g�^��{2�~��o���`����r��39[��@1��A4ة���Q9������������~J�6�ߛ�l%/�d���1������x����퇸���S?��Smkb���d�]|���4Єp��7!�[So�΍?nG��<�Eֿ�U����Z��_o�'�o�%����z��בק��1�-����s�y\� A��Ý�� �$ 䨓�ei��er������s�y��"Ꝼ�� ������y��Di��
~AxX*.d4��7l�
r�oR}Mmv�����������;9#��Y&_�I�ԫ�j<�:��u
ê/lmm2�]4
 5�:l��՝�Sg��Г���׎�D .P98#o#��r�ɭ����[?</.�|�p��ǮN#'~<��!�|$|Z���JG\R�K����Rφ�Н#����ulq�	 nb���k���wV�/�ca��2<��F�zD���,hf�ҝ�~J2#��V6V�	9��������>��^��<v5�
M
q��J�ˑ�Z��(6z��������"z5>�l4^���|6��
��Ou9�8�rO�<;���� 2��x& ��� �жWoNɵᰮY���9T��F��5�