�PNG

   IHDR         �w=�  IDATx��,G EgQݱm۶=�m�v�6�߶m�m���^*^{������w��0��O�X=ICL��%p7�s&U �a���hlcO�<w���d.�D�*�߇PG	�|Hu� ��`本QҲ���o/�n�*9��d�0�y� J	C!�e1;��5.���$T���֪ľ�ނ���s�[�/��
3�jW��5Um�#A%�6,EA����A��=���ke�E���mX�uv���y�w1���h�ￇ��9�a��y{�<�'W��pJwF���}�$��?âa�;kX�1��0��.Tɏ���{��!�>=�s�����簨�[�1�L�L�>������-a3t�w!����ލ���M�6xPM�ֺt0�ݏ�����P1b��s�`��1�g|�59D��T� ~�q#���j�Dܯ -�\?Ờ��5h�K1������M�WD���b ʿ����񠒆ˆ�JI�"�N�Rp!�{�lݓM����a�#%&��ga-x_n������-&���v�e��P~v�����W���7�;Ĵ�z}tׯ����ݢh��"2�1{�ps� �>���[����a��5�	�����դ��{.�~���Mo�)Z�b♈�|
6��M��[�+*�Ӫ��{NU}��t#ǝ�9��O��? ;���-���ӹ���'c����H�p/����O9�n�+׽�������~T��oF�w����#��0��)GS��D�<�&O)�U�(s    IEND�B`�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  <svg xmlns="http://www.w3.org/2000/svg" width="22" height="22" version="1">
 <g transform="translate(-1,-1)">
  <path style="opacity:0.2" d="M 3,2.5 C 2.446,2.5 2,2.946 2,3.5 V 21.5 C 2,22.054 2.446,22.5 3,22.5 H 14 L 22,14.5 V 3.5 C 22,2.946 21.554,2.5 21,2.5 Z"/>
  <path style="fill:#4384f1" d="M 3,2 C 2.446,2 2,2.446 2,3 V 21 C 2,21.554 2.446,22 3,22 H 14 L 22,14 V 3 C 22,2.446 21.554,2 21,2 Z"/>
  <path style="opacity:0.2" d="M 14.98,8.4996 13,8.9996 V 9.9996 L 14.992,9.4996 V 16.5 H 13 V 17.5 H 18 V 16.5 H 16 V 8.4996 Z M 7.5234,8.5016 C 7.0804,8.5098 6.7088,8.5445 6.5,8.5445 V 9.5445 C 7.0825,9.5445 8.0161,9.4352 8.7715,9.5953 9.1492,9.6753 9.4573,9.8152 9.6602,10.021 9.863,10.227 10,10.504 10,11.021 10,11.572 9.8901,11.899 9.7578,12.095 9.6255,12.292 9.4636,12.39 9.2324,12.459 8.8628,12.568 8.3365,12.512 7.8477,12.492 7.7545,12.489 7.604,12.46 7.5313,12.462 7.4624,12.465 7.404,12.468 7.3496,12.474 7.3224,12.477 7.2967,12.481 7.2637,12.488 7.2307,12.495 7.2151,12.472 7.0742,12.562 7.0566,12.573 7.012,12.607 7.0117,12.607 7.0114,12.607 6.9318,12.697 6.9316,12.697 6.9315,12.697 6.8555,12.863 6.8555,12.863 6.8554,12.863 6.8496,13.089 6.8496,13.089 6.8497,13.09 6.9276,13.271 6.9277,13.271 6.9279,13.271 7.0192,13.37 7.0195,13.371 7.0198,13.371 7.0698,13.41 7.0898,13.421 7.1099,13.433 7.1279,13.44 7.1426,13.447 7.2597,13.498 7.2778,13.488 7.3105,13.492 7.376,13.499 7.4272,13.5 7.5,13.5 7.5691,13.5 7.7451,13.48 7.834,13.486 8.0373,13.492 8.2439,13.491 8.5215,13.55 8.9086,13.632 9.304,13.786 9.5703,14.009 9.8366,14.233 10,14.495 10,14.978 10,15.478 9.8518,15.74 9.6074,15.955 9.363,16.169 8.9806,16.319 8.5332,16.402 7.6384,16.568 6.5825,16.457 6,16.457 V 17.457 C 6.4176,17.457 7.6115,17.591 8.7168,17.386 9.2695,17.284 9.8245,17.095 10.268,16.707 10.711,16.318 11,15.714 11,14.978 11,14.225 10.665,13.621 10.213,13.242 10.129,13.171 10.027,13.175 9.9375,13.117 10.167,12.983 10.42,12.9 10.586,12.654 10.86,12.247 11,11.707 11,11.021 11,10.302 10.762,9.7147 10.371,9.3179 9.9801,8.9211 9.4759,8.7222 8.9785,8.6168 8.4812,8.5114 7.9665,8.4933 7.5234,8.5015 Z"/>
  <path style="fill:#ffffff" d="M 14.98,7.9996 13,8.4996 V 9.4996 L 14.992,8.9996 V 16 H 13 V 17 H 18 V 16 H 16 V 7.9996 Z M 7.5234,8.0016 C 7.0804,8.0098 6.7088,8.0445 6.5,8.0445 V 9.0445 C 7.0825,9.0445 8.0161,8.9352 8.7715,9.0953 9.1492,9.1753 9.4573,9.3152 9.6602,9.5211 9.863,9.7269 10,10.004 10,10.521 10,11.072 9.8901,11.399 9.7578,11.595 9.6255,11.792 9.4636,11.89 9.2324,11.959 8.8628,12.068 8.3365,12.012 7.8477,11.992 7.7545,11.989 7.604,11.96 7.5313,11.962 7.4624,11.965 7.404,11.968 7.3496,11.974 7.3224,11.977 7.2967,11.981 7.2637,11.988 7.2307,11.995 7.2151,11.972 7.0742,12.062 7.0566,12.073 7.012,12.107 7.0117,12.107 7.0114,12.107 6.9318,12.197 6.9316,12.197 6.9315,12.197 6.8555,12.363 6.8555,12.363 6.8554,12.363 6.8496,12.589 6.8496,12.589 6.8497,12.59 6.9276,12.771 6.9277,12.771 6.9279,12.771 7.0192,12.87 7.0195,12.871 7.0198,12.871 7.0698,12.91 7.0898,12.921 7.1099,12.933 7.1279,12.94 7.1426,12.947 7.2597,12.998 7.2778,12.988 7.3105,12.992 7.376,12.999 7.4272,13 7.5,13 7.5691,13 7.7451,12.98 7.834,12.986 8.0373,12.992 8.2439,12.991 8.5215,13.05 8.9086,13.132 9.304,13.286 9.5703,13.509 9.8366,13.733 10,13.995 10,14.478 10,14.978 9.8518,15.24 9.6074,15.455 9.363,15.669 8.9806,15.819 8.5332,15.902 7.6384,16.068 6.5825,15.957 6,15.957 V 16.957 C 6.4176,16.957 7.6115,17.091 8.7168,16.886 9.2695,16.784 9.8245,16.595 10.268,16.207 10.711,15.818 11,15.214 11,14.478 11,13.725 10.665,13.121 10.213,12.742 10.129,12.671 10.027,12.675 9.9375,12.617 10.167,12.483 10.42,12.4 10.586,12.154 10.86,11.747 11,11.207 11,10.521 11,9.8018 10.762,9.2147 10.371,8.8179 9.9801,8.4211 9.4759,8.2222 8.9785,8.1168 8.4812,8.0114 7.9665,7.9933 7.5234,8.0015 Z"/>
  <path style="fill:#9bcdff" d="M 22,14 H 15 C 14.448,14 14,14.448 14,15 V 22 Z"/>
  <path style="opacity:0.2;fill:#ffffff" d="M 3,2 C 2.446,2 2,2.446 2,3 V 3.5 C 2,2.946 2.446,2.5 3,2.5 H 21 C 21.554,2.5 22,2.946 22,3.5 V 3 C 22,2.446 21.554,2 21,2 Z"/>
  <path style="opacity:0.2;fill:#ffffff" d="M 15,14 C 14.448,14 14,14.448 14,15 V 15.5 C 14,14.948 14.448,14.5 15,14.5 H 21.5 L 22,14 Z"/>
  <circle style="opacity:0.4" cx="6" cy="5" r="1"/>
  <circle style="opacity:0.4" cx="18" cy="5" r="1"/>
 </g>
</svg>
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �?Ў�^�6��rIY�s��R�����+nK�?z�I�w��b�2��
DS��o��4eq}������H��m-Ϧ|D	`� ��xQ4$g���J��Q��(6�R����4tsh���N�l�簄�fYL��srEk�)��:���4u.Xl����a��؇P���^�qY�}���D�K�?�N(�:��©L��uP��
k�K��r��R�<? )>Q�T�U.�YM�}��$������AL״�
:u&jj��G`�x���[8�w��� +��y�z3���P�y'S�t�8̴��c@)y觲�m���͛3.�[t�����9ĔH{y{b��f��Q��yh1�0nq#��Z] �u��%8�=J�&����'�b2�q�9��Y?�_���#��n�č�?�ܚ�p	�6tsM�siY�70�|=�w��t-'��?9� ӎ�y�l�(�TU�Y�׃��X\!ȑ�����({�h���܏��f�1������\�7G���	�oD�������pو4�p9>��k�R�?A�6�o́��> �G�,���U}���/�q�ې�Z��7���M9\�b��d8&�\���? ��N�μ�{���{q��2j��m �
+/����LN��3ma�l�y�IJQ��cI��C�X�P��r�����;�Vd�zM3�59D�{��#�,C��Z�:�.���?>�&�IQ[����="����i�"q�R@��I u)<\?;�����%�=R���cw��Ζ2�%0�}Apw24�@�O��8��V�FN���V��L�'���u=Y�ޗ�!����(�ڔ�Z�:�r�M��0�A�
��iO���(xd���-ˎs4��5p1��8����T�����6�x�U^��6 ��� ���BQ���\�C� ��j&̪�U�Nj�J8*�޸�^?p�А͸�����6Ĩ�:��;:o�����~
��	-�H��S��k�����s�L�Oh�yVi�������A�
"f
k-&|h�yu���s�z�I<HpG'Wo�K)4�Y�ܱ1$�J��}���)!�_u�����49grx�����EkP��*�G�d�W,��ո~	]�!��R$�Z�e���$�oޓ� :���|�A�<�! L��k2�mt���K��e{ Mss��F�������Ҵf�_:�V�"^qq46q�g�,��F��؇bMw)=�I���C��Ռ�Q�
���,-"B�D�z�q��y��<ΰ��b�Sq�w���Ge �j���"!Z�
@��]����D���R�[N�¿Z�O�"l������ـg.�dV	!��i�˲�K+�l�W+pg�������F����S}=�Eh�[��SP.dQKR��v]����4v�zj�#rY&��`+�z�/Z�r�{φsuRa�Ux�RG��3��+�KWIt�z� ��'�t�͎c*�\Q�7��ϔҸ3�)`T}n7)ļK���esD&��vc������im8;�0m�ul�4#��+�/����&�����*� K���bv��>�uE��A!�b���Qm.��nƟ�\R�,�eeA���,�[T0�IoE�~J�&!b`DL����w��P����-/U�4|�b>Ѯ���' ��Q�oy�Y�-	'�b�*r@C/�
�ת�ݕ�ܾ�Ԃ7�� ��	��fȻC�~]E<�,�]����+���۸�>������B��.����a�,.�5�X��h�I�� �鵭̂#}�
"���)fp��RZS�B�B{�:6=ߠ��_Z��o!��ak��rve�\�����ͼT%SA� }����b�E�UQ���ꂃ���+�J���p:�_�xp�fK1��5ʾ=��s9��F�!q��`���-��ޜ)D�BB�Q(a=�:.S�e,��@�gq���dA ��~|w����Nyᜐo@|6�JЄ����y��2Rʿil7Tm��O�����̒�k�'fw&{���� &��o�%-o�t��u����� &�T�d=�ή��+6�ȵ㣆,�?���P�H��܊����!��,�\��a�ƻ�Zv�c8�����))�/�U��~�re�yj�.D�6쉖�2a����	��y��~�L��