|�
��	cr����ܬ��پ���2�||��G��
C�$��G��=x|�����>d":mY�~�1 �����jN�!ϩJ|�p/��6r�����'�(�y,���z�w�wh���)]������n	����)nՅ[[�U�]�VV�"�b���҇��]��	�4�}��/lE���v��¼T6�tM�}��G]��I��r�3ǝ�L�U|	]�u��[-or��\���r��z�Q��o߹8�I֘ܰ���}��u�j�%��f�8vܨ���c��:�'��t����햼]<��T��u��Vw�ڑ�>RU��o}��{�f$���o����~G%���]�#؎_����_Pݹ�����n�K��k�.�����|ӕ�O
��*�j�x�֤Ĺaպ������rmʠ���?/������!�;C�PhIbB�"R�z ���Ya�,� C,"�`B�҄ T �[͛���ŷo���[}�p�J[�ݷV8a�o%u��VR���[I徕���[���޵���br��������y�1���]��
kƉ܊ni��3UJ���-����_���ʃpl����s�x�o��[MzT|d���[u��1�2�-�>��n|Ѿ ���u��n�v��ٜ��[oZG��[��@/�[�Ж�.�S5��\S��6�:}Fy�*��������!>��9�1��O�GL�8�ݶ�mN�sE��1a��9lumr��}��!�G;�U�kw�I�
˗Qw	;Q.�Z�a�L�C�%�xiPN��&(>���1��w?)M\3�i;��䎞g3����.�:�Tn��)�f�S�q�Q��7�Gnf�7�7�Zn�x��w�RlB��Cq{l#�;�Z����Dy�o��U�V��p*�Uɡl�L�����x�WK��Af�QvcW+�/�n�8iӰd��s�5�7�Pn�Q�3>������/���^��7'��:��KcP{��w[�v��h�q��P�m�5u�����xSV̙��k�s���<�b���]F��t��'���t��dP����8��!��Q{Ե(&��/�9j���
����Ow.�ȶo�JI�TV��dw�d�ȏr��f���Y��{h����v�zݎ�<������]��6Xۙ⒮fk�K���);e��b�~�'��"9�{̓��Z��i��D��s�����O��۰���?�>4����I��Js�'������c6��6��o��wT�o�"ݫc��S=��Vw5�c���WK	��D��+��BS�O:��h�����ܠ�.�D���ʎ�ُ��#/,�~4uo�3��~4�v��eqdc��7>���x�E3C�n�:��7v��[��E[�=����z�ԥL�Ǝ7��U� �������5��W<D�	�˱�d��͜�-T�V�u�7�3���y����?�f6 �ӥ��������/��^��axA,۝�~���j|A�xk�x@�>��y�bm�a����Z��{|���/���hr�;�����^��C�rD��EpV����I:i8-�|��v'��+%�v��!�ֲ�Cq.�G��C�+�wG:�V�	S���,lN�W��&�����+����=�ؒ:�CBh?�� �	R �(RF4�G�G�o��-bb��(�5t"Y����B�ȳdB����R�,��Y���ɸ��N���%�=LO�t�=]˾W��w#=���h��S���:ϙ��G�7y��	��V/z�b:��Ӌ���N/���^O/��wz9u'�Ů��%o/=y%�EHs���V�::=�3	|��ӓ��S��N_�Æ2 57�Ĺ|�&C� ���&�������zk á���Yr�)Rt�)hr�
��S|�k
��]��k�����M�k
N�5<��k�S��ҧ�R*c�z"1��;��zRzB��UEJ�9I�����t�g��d2���\"ZS^�qn"pz¹��������>�1�<��m��W�-Ū�	�<��Kt���D�(>���cߒ������'���0�7S���?��M��	����3A}F�@B��x����H��j�N (W=�pK�E��-_4�g  \�-�3��n�[P�?�<UQ&��0
���I�]$贴y�{�����~�8������x?xi�~ ����t3�9�L�yARV'L?�9�)�P�_�G,�7�t8����L�QN{�m�X���h�=����f�	��R���8f�1���~g֋a��� �o�1��%�����T���tǬ1]��cJ�r�8=���1�c#�cY���A�����g)߀����+92��p	�.�y{��O���j0k�#�.M c�%9�D!jUHx����!�s1���C"�u[�_:$�ʗ����C"WuH�7���=&d�����E=!A���Z4$R��!��� ����xøWءO$ݭ!P�6t����'���<�{�^3%�.� M��!�$���"�?����L��,�w�����qB���`*���ܾ3�c������L����7����ޜ�2M�5TW-�K���c0��3�`;��.]*�<���)��?�tZ�j���ch:�C�0�c�'��g��
8N�k������u=�	!z����TB��i�<G� �V��;i�w��:��`X��_���#�2���~�W�8�C��g�,{�Y���O ��,���Y�l�ջHpK���G`[R䭀��1C|z���vo�U��&�/#�5�ݬ�ݺ�?huw�4=���E�K���S0��%s��W�n�@�/�(�}�����mո�k�$l�g\d}[s7
�eR4��j�r۷�}}�ཛྷ����W��^-�E����+�l��n�B�`���S�ky������@Aj˩�������p�(�dC��kU��&}W9�Oe�X��;���y[T�m��L�՘3���+�<^��=�yK�y{�<����y���<o�5۽��y�0����d_��)�a�Q�&xk_I�&���0��f��T�vE;L���$��o+�n�:��I��RR�W��:;L�ov�a��{ϩ*9����w���0ux=�y��&���Tm;U����$e}}[��xk-�T�<�������3���o��o�-����9��v�tÄ���a�4��W��|��0�*��y��sa��ܨ������OUe�T&��|��[�[|}ۼƍ�0�;����y�7��

�	_y�'���i������y���}����W���v2����>�y��K��w�0ִbqTƍ�J��_�9x�����:�ZE;Ԙ��x��M�S��6s�z���J��_�M)�;���_I��R%"�.=g��U�w�ʸ�*���]M��R����3؍Yr�j'�:�*�g�l3�����b�F5���}����=P���F�>�t�;s����)O-��߳K}W�{����E���=_Ǡ����E8��_|�<a��|����*�UE�_M韃��k��O�Bp1����𑇿�����|>�4�����]��g��+�#���G|�%3�'�����[w|�'��n�?��e�s�W�]�I���2��_��.����o����#��"���H�T>Н	x��:z���̸��a�4Me_��������s����|~�7>��_�s���|��|�O����ύ��B��{��|���o�oO������.���m9�}�O�{>������5��_~̗�����c�g}�������=_�o>��|�o�/���Y��[_ ��>��.��U���*O���П}���{>������5��_~�f����	���}�g������q~��|��0?���)��_���_�g����=o�o~��|�o�/C��֞Ӿ�������_�:營�}�8����m��߾̷��c>�o�"��U'�Fٟ}�_��|Ϳ�9/�i��|���[��J}�����٧�u��o���|�O��i�o����*/�����_��|�����4��.�`�ij��                 �4�  �q��`1f��,���7� ��0І�1pd4 \0����C`xO��a���ox��?���<��rG+�<���?�I����;�T�@�i:��@Z�{@�K��q *;��+t@%'�xU8�h!�*#:&�k����-���v@Ҟ����~1�E� �/a�W��=���TX��Y.�h(a���]���u��8�����=�F$� :-��t"S���٬��"H�Jͼ���n����k̓O5x8�Ph��o�Hh��z�O6�c^�/��N�(R���ˢ�b�X��@e/��t�7=y�Z*��T�4�q�L(������� : �YK<�ґ�@fx��? ��AF}�t���Ν�b�E�Gkɖ�Y��.+��Ҕ`� �����{��.��P
� 0� ��>zD�A���A����� � ��b_�GH1�00������Ȗ��^d�]�Eߌ��c#�8~?�h��`��)iKe4u���:�&=t
X�	��g[ �� Q�]�` ���T">�\?<�n�KFS�Fz�*bĽ�þi� ��#�0p�ZJZ�.=ړ$uʢ�Z��@-��,G�&���\_�3��6��Ir< YSV�act)�T�,��e�dy�dyTH�G�4�P�}��[��*��S�t_e�A�'���tRH�f��|�#�u�P��H��^���2�����P�jz�C5�H;�ֹ3ɩ�W����@$�����|�.�n�� R3k^$����I&���V��;��q����J�U$�[ՠ������]����Q��^Y�j!�lFKC�cO�ٌw`�V�L�e+m�GSEg������=��z�u]u����,ױ̎�������Q<�&�u���uF�ѝ�P�]�e+�e��\G��^�Ϩ���8�ha�8^Nf�*�c���aC�.�q+SFm%�u�@PQ�Ms�x�����q��+0�P�)X�a<G|�(qC�TTX�Ҟ�ǜ��<�l���J�bg,��8k�_9�;�����h8����&�m���ΠM����9��6��X�}����Jq������Jg��{����98�d묱aJ�j��K9��r��<�\wԗ��T��IL�T2+㎭�>vl�c����N�Q�3�y���� ^�j����Xuf!}���ֺ�:|Y�fɓ �m� �إ�r�5X���P��(<�&+�x�4�Q��:F��-�C��)�G|L9�P�M�HV���qӎ�{������^G5�:{%9zKi�T�4�Bp���/���2�|��^�u��~�Qp8vu�cv����G�u��n�!��2�u��a��b��A˅�|������G䬼�|hhny���J�Ď�&���"R�5���"��-g�A<��%��s��J��Ǐ]��� �cF�8�����?O�ՃdOy��R8bfj<a�� ��d�;ݐ�ϱ����(��A�].߳�I)�c�Vj��8v����rX�쳖�M702�?�mx���Bhk�N0kD�1�P��j���i<x�nV
���-R2%���:v�X.|��x�Zj��l�ֲΩ���1�|��ڪ��l�cwOa�"�Q����-���)�CVj3rQ��YW��П�l����C��v4rG3���,�cZ0"�u�y�m�����E8�pj<�qE�{4���"�1���
4���=*�H���3+�̞9�b+5L���XPh%�E���G��#�2@e��<t>���Q{P�p��O����!!k�*�X��Qwl^,Ǿ�-��A<���$a��Z�Z�q��4 [i���Ql�cd�(�Q�Av�H��-�4�Ǭ*��(��܎:����~��������v#���?�R������9Ijj<���٤�Y��f���Y�?~�ΉVOM�yw�/�	�9�f��Y0!Q:��7ÊHB
��NN۠P�Ӣ�A�ax�x�Ψ��ӌ`
\.��+��)�� +o���tj��1��a��j��Ų��x�G-�:ˣ�o��g��� |��H  �Eg+:��?v��7�˖3j�|</~�Z�rF���"bœF�0t���ѱ{ُ�;"�JJ�lM�w[9+9v=r�A���R���64;a���s�����p�-�]8���Gΐ�o��Oٚ����[n
G5�f�����7FC_i�#��������cl�G��xX:��*u촎?�:�hz]��}&�E�rf3�����K�u]eQ�� ��?h�����b��'ح��!]�(�b�e�Ү݌c�������m�ͨ?�΋u3u�Ў��6�K���P��Gѱ+�f�̽��Z���16)Dz�j؏ى�^B�E^�k-��Ѩ��i,?�6u2�����6�1��ˁ���Q��Q��R�^�����hc�4�<��Zlz�e<G)��$�Cp�4vc7��c����^����:�A��#C�DMRg!�A#;)���-��A<�6���(��s�YAH��vQ+��2�;g�,��1��i�f������]臢 �:lN%8&���?f�=�a)1�9�c�Bѱ/��{cznIR�h��O��)��+*y!���HȮ�s�nE�̮ĸ3�t�m�@����:���zG5�?Bp�@�H�UG��s���c�^�3��,���aU�	�?v	��uC2Sׅ�W�O����>̋~(q��\������J`G�ʓ;��������cx6T-�d�s�.�Q9#��Lm��i�52Ok�E�,�����.`�LX6<���'�Y���c���`���IG�-���;�U�لQ�n�c���t��w��[`��:ҕv.axz�Rs-ձ�H��kHE��`���x�Ѣ��[9�A� �VSu�5�5TGYX�� 
7{�	����=����_� ���Xi�|Zy ��������N+:�1��-쾊�2s3jΈ��YB[�A[�����U�Q�����e�0��"�kp{��Mvz'�@��K>��*V�х��5��˸��P!E8{�Y��$�6r�3V@
W:�M�=�I�J̓-�^��Zy���j(���V�|��I�[0�C6jE8�*
b8�1<-[�m�*� ���ux�=U\��l����ݼ�w.��-��A<�^h�7 |��ʤCz�B�,��Zxq�-��",��3j/��Y�����_�=��km�TC��s fߌ��;J?3),�
���3��>Ǟ0�Ξ����ӟp��V�2��1eIO�DB��Νt�1�A�
T��V:i�)�~t��c�XC�
��/bDh7�(dVst�UF�����t،xc;]�O=�T�+�j��:vX��}�"i'�i�a�x �h�ӏZ.|�|��1��*%C�� t�H8�'	+�Y�⫲����M�?r3j�s���,\�!?feYZ�Ih#O����m砭E����$�U�?'{Dsǧ�%w_�9���S+	�b%��PF$BQդ���[��x��Y��M*fG�娻|w��G5���?jv���u#C�MEt���c^�sd���l�)l0fx��O\�9>����e}Z�8d��Tq�iI�@�Ż����_ˇk>��J��&� 4�E'�(�@686��,��.{�2��0F<�뇟�r.��G�A�fԪ �r4�r����i����4��h^�Ó:��ĚJ��u�I��g��i����*��e�d,w[2A�)�?Bq7��x�h�I������{��9�H���+��̌�e=���]��2��R����{�UH8��Ϭ?���4�0,��[��ؔÄaJO��b����$-��A<��°�sŷ�o�'�	�)��"���q�d�chXAr͘9���䦶����h6q d,�Z��q���cw�I�9��+@[Ჭ=�8��T�Q�Pq'<�����ej�EC~<2�pA�EXA�d0�ڊt��T�p+���P]NbI���oy��9K(���.tM�҄����tIUK׿�������]ǯO��n�b�����3�������|��_��%gb��6�6O���m^,5�����l�m�,g�^�9�+c�Jt���[f�s��g&�CV�SV��D�
e�^#�d�������������F�X�Zl	�\���i5�q�#��e��	R:�Vj�|M�\�r��V�+�2������p@���~�M���bŨ��4�]�/���(��)���Y�ծ�]����|��V.��e?���Ͽ3V��9]�b|�d�Ff9�e�;���.*:0n�$](��Q麛��.:';����£e'ml�j��#���6Y+;Bh4c�Yi��_����5z?��z2� c��h�Nx�����p�%��q� �H{-���5�o��9u�;.����]wۡ�t A(�y���r���x���K֊d!$U�r2���W����JX��)A�q;��l3�ʠʔm�[�y�˰��V  r��zV:^C,p�Uԙ�l'e)f��i��.��֭��eYX+�Q�+����g}�B��0�<n�������
�a�ʂ�^�8����]���i���.o��W��l礀*�^�U��c��
�kW�����/�@G��%l���Kɍ�<G02k?�~����f����T�
����y���3���H�]��Y���ʵ�,��3�6�m����x5�W澲�
��c#�A����Y)%���HZ$�h�/[��ޮ�|�47Z�Ö��7�QKG �Y6b�pI�i�Э����"*]iq@�п9 ޢ�5F�Hd�ȩA��y�B���N�!`��x�d�����+�-�gw#�(>d�BK Y���7ΨQ�wb�JK<