�PNG

   IHDR         �w=�  $IDATx�c�#I E{gc۶m۶m[�m۶m۶�dm���赍�s�~�\�?�����c���۞�g�82���˞��+��;+P,��n����>%�x�39�4��O�p�gv9r~��w-zL��Q�A
!Bw�g�W�p���|T��w�	>HY��@��'`�;����v��5��=���N[.�:��>�D��H���~��w��*t�J�f��R�Yu�-�6+��	ϡ(x�a���^���H/!T�Io���8����v+�f��|��̸��1��'�	�~x��!�-��!Hz�'�'�x���Ut%��U�l7�n~�֐>�b�d���)��A��RĶ8d?[��d�	�����P{���p�S~�|��-/�l�d\	� �]P��	�u�	L�ͤk߁�D����\�}�&��J������A����aEBzl�e2���A�*<���%λL�f��䛦d�5Ԫg!P�']Ga�6��{/��ZD�7��Zq�t���л��T��$��TA��/����y�u�&�.cP�K֩�/֪3k���U��\
�k�x>d�F�4��>X�n*�^�V��l�ZuV��W��3���2�!E��(z�O5Ia�"<.�n���=8�>
kTX�_-�h�p:�߲p�~ۼ�-��Z�D�6J���q/jV��s��G�Q��}#���5-9`b\�'U=g�|��`,}@gO�Jͥ(����p��F�;����k�٢t9��8B���I����ȎF~,�'�/�����`O���bX�湣�    IEND�B`�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   <svg xmlns="http://www.w3.org/2000/svg" width="22" height="22" version="1">
 <rect style="fill:#ffc543" width="20" height="16" x="-21" y="3" rx="1" ry="1" transform="scale(-1,1)"/>
 <circle style="opacity:0.2" cx="6" cy="14.5" r="3"/>
 <circle style="fill:#ff5100" cx="6" cy="14" r="3"/>
 <path style="opacity:0.2;fill:#ffffff" d="M 2,3 C 1.446,3 1,3.446 1,4 l 0,0.5 c 0,-0.554 0.446,-1 1,-1 l 18,0 c 0.554,0 1,0.446 1,1 L 21,4 C 21,3.446 20.554,3 20,3 L 2,3 Z"/>
 <path style="opacity:0.2" d="m 1,18 0,0.5 c 0,0.554 0.446,1 1,1 l 18,0 c 0.554,0 1,-0.446 1,-1 L 21,18 c 0,0.554 -0.446,1 -1,1 L 2,19 C 1.446,19 1,18.554 1,18 Z"/>
 <rect style="fill:#4d4d4d" width="16" height="4" x="3" y="5"/>
 <rect style="fill:#ff5100" width="2.625" height="2" x="6.38" y="-9" transform="matrix(0,1,-1,0,0,0)"/>
 <path style="fill:#4d4d4d" d="m 12,10 a 1,1 0 0 0 -1,1 1,1 0 0 0 1,1 1,1 0 0 0 1,-1 1,1 0 0 0 -1,-1 z"/>
 <path style="fill:#4d4d4d" d="m 15,10 a 1,1 0 0 0 -1,1 1,1 0 0 0 1,1 1,1 0 0 0 1,-1 1,1 0 0 0 -1,-1 z"/>
 <path style="fill:#4d4d4d" d="m 18,10 a 1,1 0 0 0 -1,1 1,1 0 0 0 1,1 1,1 0 0 0 1,-1 1,1 0 0 0 -1,-1 z"/>
 <path style="fill:#4d4d4d" d="m 12,13 a 1,1 0 0 0 -1,1 1,1 0 0 0 1,1 1,1 0 0 0 1,-1 1,1 0 0 0 -1,-1 z"/>
 <path style="fill:#4d4d4d" d="m 15,13 a 1,1 0 0 0 -1,1 1,1 0 0 0 1,1 1,1 0 0 0 1,-1 1,1 0 0 0 -1,-1 z"/>
 <path style="fill:#4d4d4d" d="m 18,13 a 1,1 0 0 0 -1,1 1,1 0 0 0 1,1 1,1 0 0 0 1,-1 1,1 0 0 0 -1,-1 z"/>
 <path style="fill:#4d4d4d" d="m 12,16 a 1,1 0 0 0 -1,1 1,1 0 0 0 1,1 1,1 0 0 0 1,-1 1,1 0 0 0 -1,-1 z"/>
 <path style="fill:#4d4d4d" d="m 15,16 a 1,1 0 0 0 -1,1 1,1 0 0 0 1,1 1,1 0 0 0 1,-1 1,1 0 0 0 -1,-1 z"/>
 <path style="fill:#4d4d4d" d="m 18,16 a 1,1 0 0 0 -1,1 1,1 0 0 0 1,1 1,1 0 0 0 1,-1 1,1 0 0 0 -1,-1 z"/>
</svg>
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  <svg xmlns="http://www.w3.org/2000/svg" width="24" height="24" version="1.1">
 <defs>
  <style id="current-color-scheme" type="text/css">
   .ColorScheme-Text { color:#6e6e6e; } .ColorScheme-Highlight { color:#4285f4; } .ColorScheme-NeutralText { color:#ff9800; } .ColorScheme-PositiveText { color:#4caf50; } .ColorScheme-NegativeText { color:#f44336; }
  </style>
 </defs>
 <g transform="translate(4,4)">
  <path style="fill:currentColor" class="ColorScheme-Text" d="M 8,1 A 7,7 0 0 0 1,8 7,7 0 0 0 8,15 7,7 0 0 0 15,8 7,7 0 0 0 8,1 Z M 8,4 A 2,2 0 0 1 10,6 2,2 0 0 1 8,8 2,2 0 0 1 6,6 2,2 0 0 1 8,4 Z M 8,9 C 10.5,9 12,10 12,11.5 V 12 H 4 V 11.5 C 4,10 5.5,9 8,9 Z"/>
 </g>
</svg>
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �-2����4_������`e�k�
Dڄg�	���^q8m�	�K9��'b�ցH������b�hׂKu��[k�z��5��0Iع�jK��VL=�u�S��b��Qb�^�~��߸�ۉo�v$Hh/��t�&d�(����B�H����V�=�K�D�?
�}��iҜ�\��tEk������T�p�Ș6��������A"�[&�4V |k�L�[�Þ���P��Q)g�Q>����zP�Q�`;��{�/a�'H��"�D�MI0γk9�A�������A���↝3��X�V͛ �D�E�8�R��z��#m1\|P��`S�[���vg68��{N �dҀ���zˣ*��ȁ�7��툷q+�EO��{��u������~���OlK���'v��Qr���ɓW����9pB�IKU��^�k��������ډ��k#6�k�R���9>(��v,Z��]�\6�"�V�	Hb�dٽ��+�Եղ,��,���;�<|�Ǉ�NA��{��ٞy�<9�1qY1���}>�t|� �J�"��Ore����ҨU�`����A�f	����� s��$�1		�^P�%�މA���a�춍���o ��N�=��'C�]�m��2Ō1���T߄(�]���g�Uq&X�g!������Γ���p��Y&s�'f�Vl_��wzfBQ�W	y�|K1 #�)D�c�K�/�Sm��Nv�9�ח��6�k:;v��XLj��ҺߋU��jp{������E`y]���ı���T��FڐJr�r����\Oe�><^�.=�K�ܙ\Z#5��%��z�	���P/�9�)n{�rl��pF3̶�>zU$d�\:8��7�����կ�t����Rk�S3�����7�M<�p���z�԰+���$��1;;� u�ܞT�3O�e���꧌X���c��B'��m����%`��Xk"���5�=
�0�VS	B�5a��(�l�`��^�r����*\9�����Ribݑw2+���৤��a�(�G\3hj��[�}��S��M�\4W�`W���d��(���~z�	M�p�S�#8���bΊ����@��9�@W�\pQB)z[A�}�3XT��:�M Q��jX��+��*3���_�֜��V�����3F�-��P��u1[%�\y:R
�޲#G���WiL�	X޸x`���)Cp���ũv6�}�Z��3�Y�"ĊK��tB���qi��/1Β�U�Uta�˲y��Bӄ8-b�����*h�F̺������c��B�o�\�I��t�9u����Sn]=��2d]��~!a������9#�;�롍�s(:���O�~��b��td�I�s�=��I�2�;�C�D(r*�BV~��L�o�{�/��@�L�$(�n,��dߤi��J��|
9d�E_X��f������C�ZJb�H3�ӌ?D+�:(m37�iaZ�-e���"�ٓG(�=�� r�,f;I�f�������� �]/�B��d�j�숔����������~<V%�}Rj�Yz������x7�������@��������
�����:� �Q���t��'��D���ڶ��g#n���	�q$�����n�j�m�:xȃz��E�Q�����7g8	[!��9�]eU{���)�Z#�����F�ה��5�������9��4� ��B]o�=�l3I�1:����r�]�3l䳞,trP@�;�OV��B]���Z�(���ȷd���y���0�5R�"��]��$�6tT�� ��w?�	 "dK�Q��Kϲ��!��`P�U��_�-�LD5��{����9��3�F� �SM)B"�J{l�5�p&Y��>М��i<�������Rf �'Ht�鞲�M�UYK���h�9͈��zP:,�P0�u�/c=A��M��I/(�}e�E��즴h}���˲�7"ט<\C���4I�a����r۹]=θ�r�&��!U����$�G���}Qݎo����D���rKF(�՝��5N�SD9�m�4u}=sGjw$����+��.^'E�6t��1g	c!���^�&��N2�#<C�@ۛ�'��:5�C�, ,֔�:V�����Hha��c�[�`�»db��� �s;�K�CM�8��9O�[��.�R�)��<�qb)�&H��V�
^�}�O{T��y�ЧJ�]�*ɯ1`��lޤ\d�F�;�P&w`'U9��:YWn��Bz3�� P�b�1��������]K�ȏ��8�= 1D7�������~�I��u��y$oֽ�7�� ��,U�T;X��c��8��N�}��|�D����26��>�z����>�+���%+L����I�+�A@��I���s�X!�kO��m��x��AN.�mU#����h�Տ.v��Yf���iU�����c����ts0�'ǜ�C�Kk��$���	�M��G9(��H�=�)2�U�<�-��Ъ�����u2~�W�D�9QF�"�e��Z�C��3/G�������V�������5����0�B����ж$Gj0q�+ޚ례���˔[����'��y���cB;�?h�W�����9��h����e��(���x��~7I�z����#+�Y�=�d��F��9\a)�ڦ���#L����o̘[.�м"�+5�ୃ�� Q��0��[���B5�)h���R��0�%/q.}�p/7�z�%�.&.�YSfi��/B1y�����)�a�˰/~�����Bp�N�x�3t��M-p3`B�5�p��MMlsk'�"�� �\"4�@���\n���* ���wފ�#��{�/���3��M�j�<���[��ȧ���_#�g�9=5oJ�2E!��W��:Ln�)�� 	Q��]J88qjZ�|��Q6�Y��^O�ȫ�1�W�T���v�ϊQ�%�D+���Ʉ��Yo���xr���K���W�e�~%T�Q�-N�|�<1L�OH vB���bm7F�b��	5�csƷ�"�Z�?�O^vM�֎2�~+?�vT���� Ur/�=G�l�ovc쀂��}����H<��7�	]/ɢOZ�M_�"���k��cT)�ajC��Q7uCL�CF
��'��+�'m�Oa>�]S���שc�z���;O��^q+��Jرbn�	�Mg��a;?U��	���qP�-�j�WЖC���M
F(��E������Ț�6�c�A"�i����r�z��fl���<��C�c�a����㵻L�?��2re6�:�����u��dq�q.|D�b�Z��5ap��%�Wn��� ���o�����2CH)�̵���@�'h�wDg�&�̤��`g��n������i�By{�z,��\�w����;H
����ɐ�x*�6�ۄ�9�Pp����}����#E�Z9��T@�i����kP�l;�S���y|n��xE�>�~!I���+�ã����C�d�"�|�������Vm�����UA�@�a��� �����M�Q��-D)�t�d���fUh�;4��x((��r�c���w�	���f�&A��el@�1e��U-2�[�>Ǚ�0�����=!~0�a�=u���Ut�i�]R�P�3}?�ת.��p�Əx�g���nN�Q�iN��$��y�)e	!���oCM'���vz{��]z]xw�݉ '��IX�+��6F���+b(�	{2-���C9�e��CK��}`Ask���p���y�e�A���E��N�ME�=���߯��J��|x��S��-����T �6��ܺ�"���?�O���j��r��N��m�y��-u�՝�Y�lEk2�&�mBa?�|��u��ͦߨ9��4��m�Dv�SQ�yR��׺��ȷ$�y+I�]\R��rJ� N_�[�(\���Se���N��es�5���m������=et������F^��>���I6^��,V��%"�4��8ܞA�J���WG};K�����	�0���Q�!�]8@`������=z����x_��+���=��纟{�׍ഉD[y���ϵ��$0i
����h��ݦ� #���r���O)PQ�����W��kQ������t�����������W;�>��g��+e8��@��H�ม'h������n؇a�u5.ʹ��?w8e�v�/��H3����LH��Ym?��v����r�����U[U�8'�\ET��(�a�b����s�z�Xu <9����&p^kF0�����;�K�|�rb���U=�](�' Mi<���]%�c��/�EL���x0�"�����B�!��zNn�J�Q���O�pn�5�ٮ��������e��\����*�f�I���~���9a�q9��Q�2H �":������l̶�z�؅�hP�˞������thNۅE�W��dF�f�ݍ�K �Ri�!eV[�[
�ߜ���6�)�ʸ[�������� D�x
���#`O�K�,��.�����iMmn�������~v����̚�]*��v�~F�'��7|��#�ɑ������.�UG�"��C��k`��	�r�9��0���s0���%���T7�$�	X�ʖ7��# ����4��9��W��!��H�8w��0��N�rJZ�M�b$3�uJ���e���;�o�����V�Ȉ�d�t+�O�'�ڷebL��9n)(�K���R��K�yh!KO�^�P+NU�[2{�.��Y�^��؊����ǈ���������"�Utز�$���h'�b�y$�o�-��
� 4�8���Vp��M����KC�Ajw͔
K�^�a5��f��-
�v)m����F�K3�I�����K�AP�N!�\��t��.��$:�H;����7�����7mŢ�Ѽ�h�;��}��~1U��4�Z�{��3�vWߞӚэ�c۸��J[oE�I�����J�0&�J�2��s&K�OF�T�1~N��AP R����YO}� �)|3gOܶv0�X�EC��O���"$L�B���A#�>�2'�{鷏0ujGK�u���p�<	��X+Y��R|e��\�gQ585*).�⣧
-��v'"]$)�bsn>r�i@e��H�qDn���a�@��&���I��q����w��xm]�������0�4h7�*U������'�c���ʷ?�aX�~�y�*�%{�V��ےvs�^N6l:t�4��Ƥ�m2v��k�b~0 |@��q��Ͷ��p�UV��*$_OI�D�k����Ԍ�6�J�iUZI�F5�!�0�O�u��lJ;�8�jJ�[�쯜��}3�]ZΧ>:rhg���m&��n��}�ɣR:-�(7��� f�dx;����H�V2�j�	6@F)�L 